* from MMBT5179 datasheet

.MODEL 2N5179 NPN (Is=69.28E-18 Xti=3 Eg=1.11 Vaf=100 Bf=282.1 Ne=1.177 Ise=69.28E-18 Ikf=22.03m Xtb=1.5 Br=1.176
+Nc=2 Isc=0 Ikr=0 Rc=4 Cjc=1.042p Mjc=.2468 Vjc=.75 Fc=.5 Cje=1.52p Mje=.3223 Vje=.75 Tr=1.588n
+Tf=135.6p Itf=.27 Vtf=10 Xtf=30 Rb=10)

