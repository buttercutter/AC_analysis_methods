simulator lang=spice

* 2N2222A
.MODEL 2N2222 npn
+IS=3.88184e-14 BF=929.846 NF=1.10496 VAF=16.5003
+IKF=0.019539 ISE=1.0168e-11 NE=1.94752 BR=48.4545
+NR=1.07004 VAR=40.538 IKR=0.19539 ISC=1.0168e-11
+NC=4 RB=0.1 IRB=0.1 RBM=0.1
+RE=0.0001 RC=0.426673 XTB=0.1 XTI=1
+EG=1.05 CJE=2.23677e-11 VJE=0.582701 MJE=0.63466
+TF=4.06711e-10 XTF=3.92912 VTF=17712.6 ITF=0.4334
+CJC=2.23943e-11 VJC=0.576146 MJC=0.632796 XCJC=1
+FC=0.170253 CJS=0 VJS=0.75 MJS=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
